module pll (clk, rst_n, clk_40MHz, locked);

	input clk, rst_n;
	
	output clk_40MHz;
	output locked;
	

endmodule
